`timescale 100ns/1ps

module p_block128a_opt_tb;
    parameter 
endmodule