module characterRom ( Address, pxInRow );

  input       [6:0]   Address;
  output reg  [7:0]   pxInRow;

  always @ ( Address ) begin

    case ( Address )


      7'h00: pxInRow <= 8'b11111111; /*  ********  */
      7'h01: pxInRow <= 8'b11111111; /*  ********  */
      7'h02: pxInRow <= 8'b00000011; /*  **        */
      7'h03: pxInRow <= 8'b00000011; /*  **        */
      7'h04: pxInRow <= 8'b00000011; /*  **        */
      7'h05: pxInRow <= 8'b00000011; /*  **        */
      7'h06: pxInRow <= 8'b00000011; /*  **        */
      7'h07: pxInRow <= 8'b01111111; /*  *******   */
      7'h08: pxInRow <= 8'b01111111; /*  *******   */
      7'h09: pxInRow <= 8'b00000011; /*  **        */
      7'h0A: pxInRow <= 8'b00000011; /*  **        */
      7'h0B: pxInRow <= 8'b00000011; /*  **        */
      7'h0C: pxInRow <= 8'b00000011; /*  **        */
      7'h0D: pxInRow <= 8'b00000011; /*  **        */
      7'h0E: pxInRow <= 8'b00000011; /*  **        */
      7'h0F: pxInRow <= 8'b00000011; /*  **        */


      7'h10: pxInRow <= 8'b00111100; /*    ****    */
      7'h11: pxInRow <= 8'b01111110; /*   ******   */
      7'h12: pxInRow <= 8'b11000011; /*  **    **  */
      7'h13: pxInRow <= 8'b11000011; /*  **    **  */
      7'h14: pxInRow <= 8'b11000011; /*  **    **  */
      7'h15: pxInRow <= 8'b11000011; /*  **    **  */
      7'h16: pxInRow <= 8'b11000011; /*  **    **  */
      7'h17: pxInRow <= 8'b11000011; /*  **    **  */
      7'h18: pxInRow <= 8'b11000011; /*  **    **  */
      7'h19: pxInRow <= 8'b11000011; /*  **    **  */
      7'h1A: pxInRow <= 8'b11000011; /*  **    **  */
      7'h1B: pxInRow <= 8'b11000011; /*  **    **  */
      7'h1C: pxInRow <= 8'b11010011; /*  **  * **  */
      7'h1D: pxInRow <= 8'b11100011; /*  **   ***  */
      7'h1E: pxInRow <= 8'b01111110; /*   ******   */
      7'h1F: pxInRow <= 8'b10111110; /*    **** *  */

   
      7'h20: pxInRow <= 8'b11000011; /*  **    **  */
      7'h21: pxInRow <= 8'b11000011; /*  **    **  */
      7'h22: pxInRow <= 8'b11000011; /*  **    **  */
      7'h23: pxInRow <= 8'b11000011; /*  **    **  */
      7'h24: pxInRow <= 8'b11000011; /*  **    **  */
      7'h25: pxInRow <= 8'b11000011; /*  **    **  */
      7'h26: pxInRow <= 8'b11000011; /*  **    **  */
      7'h27: pxInRow <= 8'b11111111; /*  ********  */
      7'h28: pxInRow <= 8'b11111111; /*  ********  */
      7'h29: pxInRow <= 8'b11000011; /*  **    **  */
      7'h2A: pxInRow <= 8'b11000011; /*  **    **  */
      7'h2B: pxInRow <= 8'b11000011; /*  **    **  */
      7'h2C: pxInRow <= 8'b11000011; /*  **    **  */
      7'h2D: pxInRow <= 8'b11000011; /*  **    **  */
      7'h2E: pxInRow <= 8'b11000011; /*  **    **  */
      7'h2F: pxInRow <= 8'b11000011; /*  **    **  */


      7'h30: pxInRow <= 8'b11000011; /*  **    **  */
      7'h31: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h32: pxInRow <= 8'b01100110; /*   **  **   */ 
      7'h33: pxInRow <= 8'b01100110; /*   **  **   */ 
      7'h34: pxInRow <= 8'b01100110; /*   **  **   */ 
      7'h35: pxInRow <= 8'b01100110; /*   **  **   */ 
      7'h36: pxInRow <= 8'b00111100; /*    ****    */ 
      7'h37: pxInRow <= 8'b00011000; /*     **     */
      7'h38: pxInRow <= 8'b00011000; /*     **     */
      7'h39: pxInRow <= 8'b00111100; /*    ****    */ 
      7'h3A: pxInRow <= 8'b01100110; /*   **  **   */ 
      7'h3B: pxInRow <= 8'b01100110; /*   **  **   */ 
      7'h3C: pxInRow <= 8'b01100110; /*   **  **   */ 
      7'h3D: pxInRow <= 8'b11100111; /*  ***  ***  */ 
      7'h3E: pxInRow <= 8'b11000011; /*  **    **  */
      7'h3F: pxInRow <= 8'b11000011; /*  **    **  */
 

      7'h40: pxInRow <= 8'b11000011; /*  **    **  */
      7'h41: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h42: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h43: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h44: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h45: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h46: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h47: pxInRow <= 8'b11000011; /*  **    **  */
      7'h48: pxInRow <= 8'b11000011; /*  **    **  */
      7'h49: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h4A: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h4B: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h4C: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h4D: pxInRow <= 8'b11000011; /*  **    **  */ 
      7'h4E: pxInRow <= 8'b01111110; /*   ******   */
      7'h4F: pxInRow <= 8'b00111100; /*    ****    */

      7'h50: pxInRow <= 8'b00000000; /*            */
      7'h51: pxInRow <= 8'b00000000; /*            */
      7'h52: pxInRow <= 8'b00000000; /*            */
      7'h53: pxInRow <= 8'b00000000; /*            */
      7'h54: pxInRow <= 8'b00000000; /*            */
      7'h55: pxInRow <= 8'b00000000; /*            */
      7'h56: pxInRow <= 8'b00000000; /*            */
      7'h57: pxInRow <= 8'b00000000; /*            */
      7'h58: pxInRow <= 8'b00000000; /*            */
      7'h59: pxInRow <= 8'b00000000; /*            */
      7'h5A: pxInRow <= 8'b00000000; /*            */
      7'h5B: pxInRow <= 8'b00000000; /*            */
      7'h5C: pxInRow <= 8'b00000000; /*            */
      7'h5D: pxInRow <= 8'b00000000; /*            */
      7'h5E: pxInRow <= 8'b00000000; /*            */
      7'h5F: pxInRow <= 8'b00000000; /*            */
      default: pxInRow <=8'b00000000;

    endcase
                                  
  end
  
endmodule